module cnt_width_testbench; #(
    localparam 
) (
    
);
    
endmodule 

